half_adder inst0
(
.in0	(),
.in1    (),
.sum    (),
.carry  ()
);