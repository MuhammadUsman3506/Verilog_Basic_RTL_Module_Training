full_adder full_adder_inst0
(
.in0	(),
.in1    (),
.in2    (),
.sum    (),
.carry  ()
);